`ifndef _STATE_MACHINE_VH
`define _STATE_MACHINE_VH

`define STATE_WIDTH   2
`define STATE_INIT    3'd0
`define STATE_AUTO    3'd1
`define STATE_SWITCH  3'd2
`define STATE_BIT     3'd3
`define STATE_RESET_WAIT 3'd4

`endif
