`ifndef _STATE_MACHINE_VH
`define _STATE_MACHINE_VH

`define STATE_INIT    2'd0
`define STATE_AUTO    2'd1
`define STATE_SWITCH  2'd2
`define STATE_BIT     2'd3

`endif
