`ifndef _SEVEN_SEGMENT_DISPLAY_VH
`define _SEVEN_SEGMENT_DISPLAY_VH

`define SEGMENT_A 7'b0000001
`define SEGMENT_B 7'b0000010
`define SEGMENT_C 7'b0000100
`define SEGMENT_D 7'b0001000
`define SEGMENT_E 7'b0010000
`define SEGMENT_F 7'b0100000
`define SEGMENT_G 7'b1000000

`endif
